// ============================================================================
// Copyright (c) 2016 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altera Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL/Verilog or C/C++ source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//  
//  
//                     web: http://www.terasic.com/  
//                     email: support@terasic.com
//
// ============================================================================
//Date:  Wed May 11 09:51:57 2016
// ============================================================================


module DE10_LITE_SDRAM_Nios_Test(

      ///////// Clocks /////////
      input              ADC_CLK_10,
      input              MAX10_CLK1_50,
      input              MAX10_CLK2_50,

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,

      ///////// Clock Generator I2C /////////
      output             CLK_I2C_SCL,
      inout              CLK_I2C_SDA,

      ///////// GSENSOR /////////
      output             GSENSOR_SCLK,
      inout              GSENSOR_SDO,
      inout              GSENSOR_SDI,
      input    [ 2: 1]   GSENSOR_INT,
      output             GSENSOR_CS_N,

      ///////// GPIO /////////
      inout    [35: 0]   GPIO,

      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N 

);


//=======================================================
//  REG/WIRE declarations
//=======================================================

wire ad9226_clk;
wire ad9226_otr;
wire [11:0] ad9226_d;


//=======================================================
//  Structural coding
//=======================================================


DE10_LITE_Qsys u0 
(
 .clk_clk                           (MAX10_CLK2_50),                           //                        clk.clk
 .reset_reset_n                     (1'b1),                     //                      reset.reset_n
 .altpll_0_locked_conduit_export    (),    //    altpll_0_locked_conduit.export
 .altpll_0_phasedone_conduit_export (), // altpll_0_phasedone_conduit.export
 .altpll_0_areset_conduit_export    (),     //    altpll_0_areset_conduit.export
 
 .key_external_connection_export    (KEY),    //    key_external_connection.export
 
 //SDRAM
 .clk_sdram_clk(DRAM_CLK),                    //               clk_sdram.clk
 .sdram_wire_addr(DRAM_ADDR),                 //              sdram_wire.addr
 .sdram_wire_ba(DRAM_BA),                     //                        .ba
 .sdram_wire_cas_n(DRAM_CAS_N),               //                        .cas_n
 .sdram_wire_cke(DRAM_CKE),                   //                        .cke
 .sdram_wire_cs_n(DRAM_CS_N),                 //                        .cs_n
 .sdram_wire_dq(DRAM_DQ),                     //                        .dq
 .sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),      //                        .dqm
 .sdram_wire_ras_n(DRAM_RAS_N),               //                        .ras_n
 .sdram_wire_we_n(DRAM_WE_N),                 //                        .we_n

 //ADC
 .ad9226_clk_o(ad9226_clk),
 .ad9226_d_i(ad9226_d),
 .ad9226_otr_i(ad9226_otr) 
 
 );
   
 assign ad9226_d[0] = GPIO[10];
 assign GPIO[11] = ad9226_clk;
 assign ad9226_d[2] = GPIO[12];
 assign ad9226_d[1] = GPIO[13];
 assign ad9226_d[4] = GPIO[14];
 assign ad9226_d[3] = GPIO[15];
 assign ad9226_d[6] = GPIO[16];
 assign ad9226_d[5] = GPIO[17];
 assign ad9226_d[8] = GPIO[18];
 assign ad9226_d[7] = GPIO[19];
 assign ad9226_d[10] = GPIO[20];
 assign ad9226_d[9] = GPIO[21];
 assign ad9226_otr = GPIO[22];
 assign ad9226_d[11] = GPIO[23];
   
endmodule
